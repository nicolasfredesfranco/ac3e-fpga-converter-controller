
module top();
endmodule
